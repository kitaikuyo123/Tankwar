module ROM_music(
    input clk,
    input [7:0] address,
    output reg [7:0] note
);

    always @(posedge clk)
    case(address)
        // 前奏：鼓点节奏（休止符模拟鼓点）
        0:  note <= 8'd0;     // 休止符
        1:  note <= 8'd0;
        2:  note <= 8'd0;
        3:  note <= 8'd0;
        4:  note <= 8'd0;
        5:  note <= 8'd0;
        6:  note <= 8'd0;
        7:  note <= 8'd0;
        
        // 主歌第一段："在这个风起云涌的战场上"
        8:  note <= 8'd33;    // 中音C（C4）
        9:  note <= 8'd35;    // 中音D（D4）
        10: note <= 8'd38;    // 中音E（E4）
        11: note <= 8'd40;    // 中音F（F4）
        12: note <= 8'd43;    // 中音G（G4）
        13: note <= 8'd45;    // 中音A（A4）
        14: note <= 8'd48;    // 中音B（B4）
        15: note <= 8'd51;    // 高音C（C5）
        
        16: note <= 8'd48;    // 中音B（B4）
        17: note <= 8'd45;    // 中音A（A4）
        18: note <= 8'd43;    // 中音G（G4）
        19: note <= 8'd40;    // 中音F（F4）
        20: note <= 8'd38;    // 中音E（E4）
        21: note <= 8'd35;    // 中音D（D4）
        22: note <= 8'd33;    // 中音C（C4）
        23: note <= 8'd33;    // 中音C（C4）
        
        // "暴风少年登场"
        24: note <= 8'd35;    // 中音D（D4）
        25: note <= 8'd35;    // 中音D（D4）
        26: note <= 8'd38;    // 中音E（E4）
        27: note <= 8'd38;    // 中音E（E4）
        28: note <= 8'd40;    // 中音F（F4）
        29: note <= 8'd40;    // 中音F（F4）
        30: note <= 8'd43;    // 中音G（G4）
        31: note <= 8'd43;    // 中音G（G4）
        
        // "在战胜烈火重重的咆哮声"
        32: note <= 8'd45;    // 中音A（A4）
        33: note <= 8'd45;    // 中音A（A4）
        34: note <= 8'd48;    // 中音B（B4）
        35: note <= 8'd48;    // 中音B（B4）
        36: note <= 8'd51;    // 高音C（C5）
        37: note <= 8'd51;    // 高音C（C5）
        38: note <= 8'd53;    // 高音D（D5）
        39: note <= 8'd53;    // 高音D（D5）
        
        // "喧闹整个世界"
        40: note <= 8'd55;    // 高音E（E5）
        41: note <= 8'd55;    // 高音E（E5）
        42: note <= 8'd55;    // 高音E（E5）
        43: note <= 8'd55;    // 高音E（E5）
        44: note <= 8'd53;    // 高音D（D5）
        45: note <= 8'd53;    // 高音D（D5）
        46: note <= 8'd51;    // 高音C（C5）
        47: note <= 8'd51;    // 高音C（C5）
        
        // 副歌前奏
        48: note <= 8'd48;    // 中音B（B4）
        49: note <= 8'd48;    // 中音B（B4）
        50: note <= 8'd51;    // 高音C（C5）
        51: note <= 8'd51;    // 高音C（C5）
        52: note <= 8'd53;    // 高音D（D5）
        53: note <= 8'd53;    // 高音D（D5）
        54: note <= 8'd55;    // 高音E（E5）
        55: note <= 8'd55;    // 高音E（E5）
        
        // 副歌："硝烟狂飞的讯号 机甲时代正来到"
        56: note <= 8'd58;    // 高音F#（F#5）
        57: note <= 8'd58;    // 高音F#（F#5）
        58: note <= 8'd60;    // 高音G（G5）
        59: note <= 8'd60;    // 高音G（G5）
        60: note <= 8'd63;    // 高音A（A5）
        61: note <= 8'd63;    // 高音A（A5）
        62: note <= 8'd65;    // 高音B（B5）
        63: note <= 8'd65;    // 高音B（B5）
        
        64: note <= 8'd68;    // 超高音C（C6）
        65: note <= 8'd68;    // 超高音C（C6）
        66: note <= 8'd68;    // 超高音C（C6）
        67: note <= 8'd68;    // 超高音C（C6）
        68: note <= 8'd65;    // 高音B（B5）
        69: note <= 8'd65;    // 高音B（B5）
        70: note <= 8'd63;    // 高音A（A5）
        71: note <= 8'd63;    // 高音A（A5）
        
        // "热血逆流而上 战车在发烫 勇士也势不可挡"
        72: note <= 8'd60;    // 高音G（G5）
        73: note <= 8'd60;    // 高音G（G5）
        74: note <= 8'd60;    // 高音G（G5）
        75: note <= 8'd60;    // 高音G（G5）
        76: note <= 8'd58;    // 高音F#（F#5）
        77: note <= 8'd58;    // 高音F#（F#5）
        78: note <= 8'd55;    // 高音E（E5）
        79: note <= 8'd55;    // 高音E（E5）
        
        80: note <= 8'd53;    // 高音D（D5）
        81: note <= 8'd53;    // 高音D（D5）
        82: note <= 8'd51;    // 高音C（C5）
        83: note <= 8'd51;    // 高音C（C5）
        84: note <= 8'd48;    // 中音B（B4）
        85: note <= 8'd48;    // 中音B（B4）
        86: note <= 8'd45;    // 中音A（A4）
        87: note <= 8'd45;    // 中音A（A4）
        
        // 间奏（鼓点+旋律）
        88: note <= 8'd0;     // 休止符（鼓点）
        89: note <= 8'd0;
        90: note <= 8'd0;
        91: note <= 8'd0;
        92: note <= 8'd33;    // 中音C（C4）
        93: note <= 8'd38;    // 中音E（E4）
        94: note <= 8'd43;    // 中音G（G4）
        95: note <= 8'd51;    // 高音C（C5）
        
        96: note <= 8'd0;     // 休止符
        97: note <= 8'd0;
        98: note <= 8'd0;
        99: note <= 8'd0;
        100: note <= 8'd51;   // 高音C（C5）
        101: note <= 8'd48;   // 中音B（B4）
        102: note <= 8'd45;   // 中音A（A4）
        103: note <= 8'd43;   // 中音G（G4）
        
        // 第二段主歌（简化处理，重复部分略）
        104: note <= 8'd33;   // 中音C（C4）
        105: note <= 8'd35;   // 中音D（D4）
        106: note <= 8'd38;   // 中音E（E4）
        107: note <= 8'd40;   // 中音F（F4）
        108: note <= 8'd43;   // 中音G（G4）
        109: note <= 8'd45;   // 中音A（A4）
        110: note <= 8'd48;   // 中音B（B4）
        111: note <= 8'd51;   // 高音C（C5）
        
        112: note <= 8'd48;   // 中音B（B4）
        113: note <= 8'd45;   // 中音A（A4）
        114: note <= 8'd43;   // 中音G（G4）
        115: note <= 8'd40;   // 中音F（F4）
        116: note <= 8'd38;   // 中音E（E4）
        117: note <= 8'd35;   // 中音D（D4）
        118: note <= 8'd33;   // 中音C（C4）
        119: note <= 8'd33;   // 中音C（C4）
        
        // 副歌重复（升高八度）
        120: note <= 8'd66;   // 超高音C（C6，原C5升高八度）
        121: note <= 8'd66;   // 超高音C（C6）
        122: note <= 8'd68;   // 超高音D（D6）
        123: note <= 8'd68;   // 超高音D（D6）
        124: note <= 8'd70;   // 超高音E（E6）
        125: note <= 8'd70;   // 超高音E（E6）
        126: note <= 8'd73;   // 超高音F#（F#6）
        127: note <= 8'd73;   // 超高音F#（F#6）
        
        // 尾声
        128: note <= 8'd75;   // 超高音G（G6）
        129: note <= 8'd75;   // 超高音G（G6）
        130: note <= 8'd75;   // 超高音G（G6）
        131: note <= 8'd75;   // 超高音G（G6）
        132: note <= 8'd73;   // 超高音F#（F#6）
        133: note <= 8'd73;   // 超高音F#（F#6）
        134: note <= 8'd70;   // 超高音E（E6）
        135: note <= 8'd70;   // 超高音E（E6）
        
        136: note <= 8'd68;   // 超高音D（D6）
        137: note <= 8'd68;   // 超高音D（D6）
        138: note <= 8'd66;   // 超高音C（C6）
        139: note <= 8'd66;   // 超高音C（C6）
        140: note <= 8'd63;   // 高音A（A5）
        141: note <= 8'd63;   // 高音A（A5）
        142: note <= 8'd60;   // 高音G（G5）
        143: note <= 8'd60;   // 高音G（G5）
        
        // 渐弱收尾
        144: note <= 8'd58;   // 高音F#（F#5）
        145: note <= 8'd58;   // 高音F#（F#5）
        146: note <= 8'd55;   // 高音E（E5）
        147: note <= 8'd55;   // 高音E（E5）
        148: note <= 8'd53;   // 高音D（D5）
        149: note <= 8'd53;   // 高音D（D5）
        150: note <= 8'd51;   // 高音C（C5）
        151: note <= 8'd51;   // 高音C（C5）
        
        152: note <= 8'd48;   // 中音B（B4）
        153: note <= 8'd48;   // 中音B（B4）
        154: note <= 8'd45;   // 中音A（A4）
        155: note <= 8'd45;   // 中音A（A4）
        156: note <= 8'd43;   // 中音G（G4）
        157: note <= 8'd43;   // 中音G（G4）
        158: note <= 8'd40;   // 中音F（F4）
        159: note <= 8'd40;   // 中音F（F4）
        
        // 结尾休止符
        160: note <= 8'd0;
        161: note <= 8'd0;
        162: note <= 8'd0;
        163: note <= 8'd0;
        164: note <= 8'd0;
        165: note <= 8'd0;
        166: note <= 8'd0;
        167: note <= 8'd0;
        
        168: note <= 8'd0;
        169: note <= 8'd0;
        170: note <= 8'd0;
        171: note <= 8'd0;
        172: note <= 8'd0;
        173: note <= 8'd0;
        174: note <= 8'd0;
        175: note <= 8'd0;
        
        // 扩展预留（176-255）
        default: note <= 8'd0;
    endcase
endmodule